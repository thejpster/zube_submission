VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO zube_wrapped_project
  CLASS BLOCK ;
  FOREIGN zube_wrapped_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 20.330 296.000 20.610 300.000 ;
=======
        RECT 19.410 296.000 19.690 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.720 300.000 1.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 62.600 300.000 63.200 ;
=======
        RECT 296.000 64.640 300.000 65.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 68.720 300.000 69.320 ;
=======
        RECT 296.000 70.760 300.000 71.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 74.840 300.000 75.440 ;
=======
        RECT 296.000 77.560 300.000 78.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 80.960 300.000 81.560 ;
=======
        RECT 296.000 83.680 300.000 84.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 87.080 300.000 87.680 ;
=======
        RECT 296.000 90.480 300.000 91.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 93.200 300.000 93.800 ;
=======
        RECT 296.000 96.600 300.000 97.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 99.320 300.000 99.920 ;
=======
        RECT 296.000 103.400 300.000 104.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 106.120 300.000 106.720 ;
=======
        RECT 296.000 109.520 300.000 110.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 112.240 300.000 112.840 ;
=======
        RECT 296.000 116.320 300.000 116.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 118.360 300.000 118.960 ;
=======
        RECT 296.000 122.440 300.000 123.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.840 300.000 7.440 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 124.480 300.000 125.080 ;
=======
        RECT 296.000 129.240 300.000 129.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 130.600 300.000 131.200 ;
=======
        RECT 296.000 135.360 300.000 135.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 136.720 300.000 137.320 ;
=======
        RECT 296.000 141.480 300.000 142.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 142.840 300.000 143.440 ;
=======
        RECT 296.000 148.280 300.000 148.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 148.960 300.000 149.560 ;
=======
        RECT 296.000 154.400 300.000 155.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 155.760 300.000 156.360 ;
=======
        RECT 296.000 161.200 300.000 161.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 161.880 300.000 162.480 ;
=======
        RECT 296.000 167.320 300.000 167.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 168.000 300.000 168.600 ;
=======
        RECT 296.000 174.120 300.000 174.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 174.120 300.000 174.720 ;
=======
        RECT 296.000 180.240 300.000 180.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 180.240 300.000 180.840 ;
=======
        RECT 296.000 187.040 300.000 187.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 12.960 300.000 13.560 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 186.360 300.000 186.960 ;
=======
        RECT 296.000 193.160 300.000 193.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 192.480 300.000 193.080 ;
=======
        RECT 296.000 199.280 300.000 199.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 198.600 300.000 199.200 ;
=======
        RECT 296.000 206.080 300.000 206.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 205.400 300.000 206.000 ;
=======
        RECT 296.000 212.200 300.000 212.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 211.520 300.000 212.120 ;
=======
        RECT 296.000 219.000 300.000 219.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 217.640 300.000 218.240 ;
=======
        RECT 296.000 225.120 300.000 225.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 223.760 300.000 224.360 ;
=======
        RECT 296.000 231.920 300.000 232.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 229.880 300.000 230.480 ;
=======
        RECT 296.000 238.040 300.000 238.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 19.080 300.000 19.680 ;
=======
        RECT 296.000 19.760 300.000 20.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 25.200 300.000 25.800 ;
=======
        RECT 296.000 25.880 300.000 26.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 31.320 300.000 31.920 ;
=======
        RECT 296.000 32.680 300.000 33.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 37.440 300.000 38.040 ;
=======
        RECT 296.000 38.800 300.000 39.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 43.560 300.000 44.160 ;
=======
        RECT 296.000 45.600 300.000 46.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 49.680 300.000 50.280 ;
=======
        RECT 296.000 51.720 300.000 52.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 56.480 300.000 57.080 ;
=======
        RECT 296.000 58.520 300.000 59.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.800 300.000 5.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 66.680 300.000 67.280 ;
=======
        RECT 296.000 68.720 300.000 69.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 72.800 300.000 73.400 ;
=======
        RECT 296.000 75.520 300.000 76.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 78.920 300.000 79.520 ;
=======
        RECT 296.000 81.640 300.000 82.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 85.040 300.000 85.640 ;
=======
        RECT 296.000 88.440 300.000 89.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 91.160 300.000 91.760 ;
=======
        RECT 296.000 94.560 300.000 95.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 97.280 300.000 97.880 ;
=======
        RECT 296.000 101.360 300.000 101.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 104.080 300.000 104.680 ;
=======
        RECT 296.000 107.480 300.000 108.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 110.200 300.000 110.800 ;
=======
        RECT 296.000 113.600 300.000 114.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 116.320 300.000 116.920 ;
=======
        RECT 296.000 120.400 300.000 121.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 122.440 300.000 123.040 ;
=======
        RECT 296.000 126.520 300.000 127.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 128.560 300.000 129.160 ;
=======
        RECT 296.000 133.320 300.000 133.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 134.680 300.000 135.280 ;
=======
        RECT 296.000 139.440 300.000 140.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 140.800 300.000 141.400 ;
=======
        RECT 296.000 146.240 300.000 146.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 146.920 300.000 147.520 ;
=======
        RECT 296.000 152.360 300.000 152.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 153.720 300.000 154.320 ;
=======
        RECT 296.000 159.160 300.000 159.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 159.840 300.000 160.440 ;
=======
        RECT 296.000 165.280 300.000 165.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 165.960 300.000 166.560 ;
=======
        RECT 296.000 172.080 300.000 172.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 172.080 300.000 172.680 ;
=======
        RECT 296.000 178.200 300.000 178.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 178.200 300.000 178.800 ;
=======
        RECT 296.000 184.320 300.000 184.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 184.320 300.000 184.920 ;
=======
        RECT 296.000 191.120 300.000 191.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 17.040 300.000 17.640 ;
=======
        RECT 296.000 17.720 300.000 18.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 190.440 300.000 191.040 ;
=======
        RECT 296.000 197.240 300.000 197.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 196.560 300.000 197.160 ;
=======
        RECT 296.000 204.040 300.000 204.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 203.360 300.000 203.960 ;
=======
        RECT 296.000 210.160 300.000 210.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 209.480 300.000 210.080 ;
=======
        RECT 296.000 216.960 300.000 217.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 215.600 300.000 216.200 ;
=======
        RECT 296.000 223.080 300.000 223.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 221.720 300.000 222.320 ;
=======
        RECT 296.000 229.880 300.000 230.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 227.840 300.000 228.440 ;
=======
        RECT 296.000 236.000 300.000 236.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 233.960 300.000 234.560 ;
=======
        RECT 296.000 242.120 300.000 242.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 23.160 300.000 23.760 ;
=======
        RECT 296.000 23.840 300.000 24.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 29.280 300.000 29.880 ;
=======
        RECT 296.000 30.640 300.000 31.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 35.400 300.000 36.000 ;
=======
        RECT 296.000 36.760 300.000 37.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 41.520 300.000 42.120 ;
=======
        RECT 296.000 43.560 300.000 44.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 47.640 300.000 48.240 ;
=======
        RECT 296.000 49.680 300.000 50.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 54.440 300.000 55.040 ;
=======
        RECT 296.000 55.800 300.000 56.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 60.560 300.000 61.160 ;
=======
        RECT 296.000 62.600 300.000 63.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.760 300.000 3.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 64.640 300.000 65.240 ;
=======
        RECT 296.000 66.680 300.000 67.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 70.760 300.000 71.360 ;
=======
        RECT 296.000 73.480 300.000 74.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 76.880 300.000 77.480 ;
=======
        RECT 296.000 79.600 300.000 80.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 83.000 300.000 83.600 ;
=======
        RECT 296.000 86.400 300.000 87.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 89.120 300.000 89.720 ;
=======
        RECT 296.000 92.520 300.000 93.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 95.240 300.000 95.840 ;
=======
        RECT 296.000 98.640 300.000 99.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 102.040 300.000 102.640 ;
=======
        RECT 296.000 105.440 300.000 106.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 108.160 300.000 108.760 ;
=======
        RECT 296.000 111.560 300.000 112.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 114.280 300.000 114.880 ;
=======
        RECT 296.000 118.360 300.000 118.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 120.400 300.000 121.000 ;
=======
        RECT 296.000 124.480 300.000 125.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.880 300.000 9.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 126.520 300.000 127.120 ;
=======
        RECT 296.000 131.280 300.000 131.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 132.640 300.000 133.240 ;
=======
        RECT 296.000 137.400 300.000 138.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 138.760 300.000 139.360 ;
=======
        RECT 296.000 144.200 300.000 144.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 144.880 300.000 145.480 ;
=======
        RECT 296.000 150.320 300.000 150.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 151.680 300.000 152.280 ;
=======
        RECT 296.000 156.440 300.000 157.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 157.800 300.000 158.400 ;
=======
        RECT 296.000 163.240 300.000 163.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 163.920 300.000 164.520 ;
=======
        RECT 296.000 169.360 300.000 169.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 170.040 300.000 170.640 ;
=======
        RECT 296.000 176.160 300.000 176.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 176.160 300.000 176.760 ;
=======
        RECT 296.000 182.280 300.000 182.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 182.280 300.000 182.880 ;
=======
        RECT 296.000 189.080 300.000 189.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 15.000 300.000 15.600 ;
=======
        RECT 296.000 15.680 300.000 16.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 188.400 300.000 189.000 ;
=======
        RECT 296.000 195.200 300.000 195.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 194.520 300.000 195.120 ;
=======
        RECT 296.000 202.000 300.000 202.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 201.320 300.000 201.920 ;
=======
        RECT 296.000 208.120 300.000 208.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 207.440 300.000 208.040 ;
=======
        RECT 296.000 214.920 300.000 215.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 213.560 300.000 214.160 ;
=======
        RECT 296.000 221.040 300.000 221.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 219.680 300.000 220.280 ;
=======
        RECT 296.000 227.160 300.000 227.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 225.800 300.000 226.400 ;
=======
        RECT 296.000 233.960 300.000 234.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 231.920 300.000 232.520 ;
=======
        RECT 296.000 240.080 300.000 240.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 21.120 300.000 21.720 ;
=======
        RECT 296.000 21.800 300.000 22.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 27.240 300.000 27.840 ;
=======
        RECT 296.000 27.920 300.000 28.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 33.360 300.000 33.960 ;
=======
        RECT 296.000 34.720 300.000 35.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 39.480 300.000 40.080 ;
=======
        RECT 296.000 40.840 300.000 41.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 45.600 300.000 46.200 ;
=======
        RECT 296.000 47.640 300.000 48.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 52.400 300.000 53.000 ;
=======
        RECT 296.000 53.760 300.000 54.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 58.520 300.000 59.120 ;
=======
        RECT 296.000 60.560 300.000 61.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 236.000 300.000 236.600 ;
=======
        RECT 0.000 176.840 4.000 177.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
=======
      LAYER met2 ;
        RECT 247.110 296.000 247.390 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
=======
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
=======
      LAYER met2 ;
        RECT 250.330 296.000 250.610 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
=======
      LAYER met3 ;
        RECT 296.000 267.960 300.000 268.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 259.990 296.000 260.270 300.000 ;
=======
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 229.200 4.000 229.800 ;
=======
        RECT 0.000 236.680 4.000 237.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
=======
      LAYER met2 ;
        RECT 256.310 296.000 256.590 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 269.650 296.000 269.930 300.000 ;
=======
        RECT 137.630 0.000 137.910 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 273.400 300.000 274.000 ;
=======
        RECT 0.000 247.560 4.000 248.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
=======
      LAYER met2 ;
        RECT 268.270 296.000 268.550 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
=======
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
=======
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 257.760 4.000 258.360 ;
=======
        RECT 0.000 258.440 4.000 259.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 279.520 300.000 280.120 ;
=======
      LAYER met2 ;
        RECT 277.010 296.000 277.290 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 283.600 300.000 284.200 ;
=======
        RECT 0.000 269.320 4.000 269.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 224.570 0.000 224.850 4.000 ;
=======
        RECT 197.890 0.000 198.170 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 282.070 296.000 282.350 300.000 ;
=======
      LAYER met3 ;
        RECT 296.000 291.760 300.000 292.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 285.290 296.000 285.570 300.000 ;
=======
        RECT 221.810 0.000 222.090 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 288.510 296.000 288.790 300.000 ;
=======
        RECT 245.730 0.000 246.010 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 258.150 0.000 258.430 4.000 ;
=======
        RECT 257.690 0.000 257.970 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
=======
      LAYER met3 ;
        RECT 296.000 295.840 300.000 296.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 241.130 296.000 241.410 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 293.800 300.000 294.400 ;
=======
        RECT 296.000 297.880 300.000 298.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
=======
      LAYER met2 ;
        RECT 294.950 296.000 295.230 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 41.490 0.000 41.770 4.000 ;
=======
        RECT 41.950 0.000 42.230 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 58.050 0.000 58.330 4.000 ;
=======
        RECT 232.390 296.000 232.670 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 244.350 296.000 244.630 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 247.570 296.000 247.850 300.000 ;
=======
      LAYER met3 ;
        RECT 296.000 255.040 300.000 255.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 74.610 0.000 74.890 4.000 ;
=======
        RECT 241.130 296.000 241.410 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
=======
      LAYER met2 ;
        RECT 244.350 296.000 244.630 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 254.010 296.000 254.290 300.000 ;
=======
        RECT 125.670 0.000 125.950 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
=======
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 257.080 300.000 257.680 ;
=======
        RECT 296.000 263.880 300.000 264.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 209.480 4.000 210.080 ;
=======
        RECT 0.000 220.360 4.000 220.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 259.120 300.000 259.720 ;
=======
        RECT 0.000 231.240 4.000 231.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 224.440 4.000 225.040 ;
=======
        RECT 296.000 270.000 300.000 270.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 174.890 0.000 175.170 4.000 ;
=======
        RECT 253.090 296.000 253.370 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 265.240 300.000 265.840 ;
=======
        RECT 296.000 278.840 300.000 279.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 263.210 296.000 263.490 300.000 ;
=======
        RECT 259.070 296.000 259.350 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 269.320 300.000 269.920 ;
=======
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 275.440 300.000 276.040 ;
=======
      LAYER met2 ;
        RECT 265.050 296.000 265.330 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
=======
      LAYER met2 ;
        RECT 271.030 296.000 271.310 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 156.440 4.000 157.040 ;
=======
        RECT 0.000 187.720 4.000 188.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 191.450 0.000 191.730 4.000 ;
=======
        RECT 185.930 0.000 186.210 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 276.090 296.000 276.370 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 263.200 4.000 263.800 ;
=======
        RECT 296.000 284.960 300.000 285.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 267.960 4.000 268.560 ;
=======
        RECT 296.000 289.720 300.000 290.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 278.850 296.000 279.130 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 287.680 300.000 288.280 ;
=======
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
=======
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 291.730 296.000 292.010 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
=======
      LAYER met2 ;
        RECT 282.990 296.000 283.270 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 294.950 296.000 295.230 300.000 ;
=======
        RECT 269.650 0.000 269.930 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 242.120 300.000 242.720 ;
=======
        RECT 296.000 246.880 300.000 247.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 295.840 300.000 296.440 ;
=======
      LAYER met2 ;
        RECT 292.190 296.000 292.470 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 297.880 300.000 298.480 ;
=======
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 244.160 300.000 244.760 ;
=======
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 246.200 300.000 246.800 ;
=======
        RECT 296.000 250.960 300.000 251.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
=======
      LAYER met2 ;
        RECT 238.370 296.000 238.650 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 253.000 300.000 253.600 ;
=======
        RECT 296.000 257.760 300.000 258.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 91.630 0.000 91.910 4.000 ;
=======
        RECT 77.830 0.000 78.110 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 108.190 0.000 108.470 4.000 ;
=======
        RECT 101.750 0.000 102.030 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
=======
      LAYER met3 ;
        RECT 296.000 259.800 300.000 260.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 24.930 0.000 25.210 4.000 ;
=======
        RECT 6.070 0.000 6.350 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 204.720 4.000 205.320 ;
=======
        RECT 0.000 209.480 4.000 210.080 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 256.770 296.000 257.050 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 219.680 4.000 220.280 ;
=======
        RECT 296.000 265.920 300.000 266.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 261.160 300.000 261.760 ;
=======
        RECT 296.000 272.720 300.000 273.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 263.200 300.000 263.800 ;
=======
        RECT 296.000 276.800 300.000 277.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 267.280 300.000 267.880 ;
=======
        RECT 296.000 280.880 300.000 281.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 266.430 296.000 266.710 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 271.360 300.000 271.960 ;
=======
      LAYER met2 ;
        RECT 262.290 296.000 262.570 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 277.480 300.000 278.080 ;
=======
        RECT 296.000 282.920 300.000 283.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
=======
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 240.080 300.000 240.680 ;
=======
        RECT 0.000 193.160 4.000 193.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met2 ;
        RECT 272.870 296.000 273.150 300.000 ;
=======
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 208.010 0.000 208.290 4.000 ;
=======
        RECT 274.250 296.000 274.530 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 281.560 300.000 282.160 ;
=======
        RECT 296.000 287.680 300.000 288.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 285.640 300.000 286.240 ;
=======
      LAYER met2 ;
        RECT 280.230 296.000 280.510 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 272.720 4.000 273.320 ;
=======
        RECT 0.000 280.200 4.000 280.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 277.480 4.000 278.080 ;
=======
        RECT 296.000 293.800 300.000 294.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
=======
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 287.000 4.000 287.600 ;
=======
        RECT 0.000 296.520 4.000 297.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 289.720 300.000 290.320 ;
=======
      LAYER met2 ;
        RECT 286.210 296.000 286.490 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 291.760 300.000 292.360 ;
=======
      LAYER met2 ;
        RECT 288.970 296.000 289.250 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 165.960 4.000 166.560 ;
=======
        RECT 296.000 248.920 300.000 249.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 298.170 296.000 298.450 300.000 ;
=======
        RECT 281.610 0.000 281.890 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 291.270 0.000 291.550 4.000 ;
=======
        RECT 298.170 296.000 298.450 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
=======
      LAYER met2 ;
        RECT 229.170 296.000 229.450 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
=======
      LAYER met2 ;
        RECT 235.150 296.000 235.430 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 296.000 250.960 300.000 251.560 ;
=======
        RECT 296.000 253.000 300.000 253.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 296.000 255.040 300.000 255.640 ;
=======
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
=======
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 250.790 296.000 251.070 300.000 ;
=======
        RECT 113.710 0.000 113.990 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 195.200 4.000 195.800 ;
=======
        RECT 296.000 261.840 300.000 262.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END la1_oenb[9]
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
<<<<<<< HEAD
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 296.000 238.190 300.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
=======
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 296.000 226.690 300.000 ;
    END
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
<<<<<<< HEAD
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
=======
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 296.000 1.750 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 296.000 4.510 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 17.110 296.000 17.390 300.000 ;
=======
        RECT 16.190 296.000 16.470 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 35.970 296.000 36.250 300.000 ;
=======
        RECT 34.130 296.000 34.410 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 67.710 296.000 67.990 300.000 ;
=======
        RECT 64.030 296.000 64.310 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 70.470 296.000 70.750 300.000 ;
=======
        RECT 67.250 296.000 67.530 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 73.690 296.000 73.970 300.000 ;
=======
        RECT 70.010 296.000 70.290 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 76.910 296.000 77.190 300.000 ;
=======
        RECT 73.230 296.000 73.510 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 80.130 296.000 80.410 300.000 ;
=======
        RECT 76.450 296.000 76.730 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 83.350 296.000 83.630 300.000 ;
=======
        RECT 79.210 296.000 79.490 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 86.570 296.000 86.850 300.000 ;
=======
        RECT 82.430 296.000 82.710 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 89.790 296.000 90.070 300.000 ;
=======
        RECT 85.190 296.000 85.470 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 93.010 296.000 93.290 300.000 ;
=======
        RECT 88.410 296.000 88.690 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 95.770 296.000 96.050 300.000 ;
=======
        RECT 91.170 296.000 91.450 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 39.190 296.000 39.470 300.000 ;
=======
        RECT 37.350 296.000 37.630 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 98.990 296.000 99.270 300.000 ;
=======
        RECT 94.390 296.000 94.670 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 102.210 296.000 102.490 300.000 ;
=======
        RECT 97.150 296.000 97.430 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 105.430 296.000 105.710 300.000 ;
=======
        RECT 100.370 296.000 100.650 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 108.650 296.000 108.930 300.000 ;
=======
        RECT 103.130 296.000 103.410 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 111.870 296.000 112.150 300.000 ;
=======
        RECT 106.350 296.000 106.630 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 115.090 296.000 115.370 300.000 ;
=======
        RECT 109.110 296.000 109.390 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 117.850 296.000 118.130 300.000 ;
=======
        RECT 112.330 296.000 112.610 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 121.070 296.000 121.350 300.000 ;
=======
        RECT 115.090 296.000 115.370 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 124.290 296.000 124.570 300.000 ;
=======
        RECT 118.310 296.000 118.590 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 127.510 296.000 127.790 300.000 ;
=======
        RECT 121.070 296.000 121.350 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 42.410 296.000 42.690 300.000 ;
=======
        RECT 40.110 296.000 40.390 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 130.730 296.000 131.010 300.000 ;
=======
        RECT 124.290 296.000 124.570 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 133.950 296.000 134.230 300.000 ;
=======
        RECT 127.050 296.000 127.330 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 45.630 296.000 45.910 300.000 ;
=======
        RECT 43.330 296.000 43.610 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 48.390 296.000 48.670 300.000 ;
=======
        RECT 46.090 296.000 46.370 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 51.610 296.000 51.890 300.000 ;
=======
        RECT 49.310 296.000 49.590 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 54.830 296.000 55.110 300.000 ;
=======
        RECT 52.070 296.000 52.350 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 58.050 296.000 58.330 300.000 ;
=======
        RECT 55.290 296.000 55.570 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 61.270 296.000 61.550 300.000 ;
=======
        RECT 58.050 296.000 58.330 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 64.490 296.000 64.770 300.000 ;
=======
        RECT 61.270 296.000 61.550 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 10.670 296.000 10.950 300.000 ;
=======
        RECT 10.210 296.000 10.490 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 137.170 296.000 137.450 300.000 ;
=======
        RECT 130.270 296.000 130.550 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 168.450 296.000 168.730 300.000 ;
=======
        RECT 160.170 296.000 160.450 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 171.670 296.000 171.950 300.000 ;
=======
        RECT 163.390 296.000 163.670 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 174.890 296.000 175.170 300.000 ;
=======
        RECT 166.150 296.000 166.430 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 178.110 296.000 178.390 300.000 ;
=======
        RECT 169.370 296.000 169.650 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 181.330 296.000 181.610 300.000 ;
=======
        RECT 172.130 296.000 172.410 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 184.550 296.000 184.830 300.000 ;
=======
        RECT 175.350 296.000 175.630 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 187.310 296.000 187.590 300.000 ;
=======
        RECT 178.110 296.000 178.390 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 190.530 296.000 190.810 300.000 ;
=======
        RECT 181.330 296.000 181.610 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 193.750 296.000 194.030 300.000 ;
=======
        RECT 184.090 296.000 184.370 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 196.970 296.000 197.250 300.000 ;
=======
        RECT 187.310 296.000 187.590 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 139.930 296.000 140.210 300.000 ;
=======
        RECT 133.030 296.000 133.310 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 200.190 296.000 200.470 300.000 ;
=======
        RECT 190.070 296.000 190.350 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 203.410 296.000 203.690 300.000 ;
=======
        RECT 193.290 296.000 193.570 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 206.630 296.000 206.910 300.000 ;
=======
        RECT 196.050 296.000 196.330 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 209.390 296.000 209.670 300.000 ;
=======
        RECT 199.270 296.000 199.550 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 212.610 296.000 212.890 300.000 ;
=======
        RECT 202.030 296.000 202.310 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 215.830 296.000 216.110 300.000 ;
=======
        RECT 205.250 296.000 205.530 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 219.050 296.000 219.330 300.000 ;
=======
        RECT 208.010 296.000 208.290 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 222.270 296.000 222.550 300.000 ;
=======
        RECT 211.230 296.000 211.510 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 225.490 296.000 225.770 300.000 ;
=======
        RECT 213.990 296.000 214.270 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 228.710 296.000 228.990 300.000 ;
=======
        RECT 217.210 296.000 217.490 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 143.150 296.000 143.430 300.000 ;
=======
        RECT 136.250 296.000 136.530 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 231.930 296.000 232.210 300.000 ;
=======
        RECT 219.970 296.000 220.250 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 234.690 296.000 234.970 300.000 ;
=======
        RECT 223.190 296.000 223.470 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 146.370 296.000 146.650 300.000 ;
=======
        RECT 139.010 296.000 139.290 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 149.590 296.000 149.870 300.000 ;
=======
        RECT 142.230 296.000 142.510 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 152.810 296.000 153.090 300.000 ;
=======
        RECT 144.990 296.000 145.270 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 156.030 296.000 156.310 300.000 ;
=======
        RECT 148.210 296.000 148.490 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 159.250 296.000 159.530 300.000 ;
=======
        RECT 151.430 296.000 151.710 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 162.470 296.000 162.750 300.000 ;
=======
        RECT 154.190 296.000 154.470 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 165.230 296.000 165.510 300.000 ;
=======
        RECT 157.410 296.000 157.690 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 2.080 4.000 2.680 ;
=======
        RECT 0.000 2.760 4.000 3.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 50.360 4.000 50.960 ;
=======
        RECT 0.000 57.160 4.000 57.760 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 55.120 4.000 55.720 ;
=======
        RECT 0.000 62.600 4.000 63.200 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 59.880 4.000 60.480 ;
=======
        RECT 0.000 68.040 4.000 68.640 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 69.400 4.000 70.000 ;
=======
        RECT 0.000 78.920 4.000 79.520 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 74.160 4.000 74.760 ;
=======
        RECT 0.000 84.360 4.000 84.960 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 78.920 4.000 79.520 ;
=======
        RECT 0.000 89.800 4.000 90.400 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 83.680 4.000 84.280 ;
=======
        RECT 0.000 95.240 4.000 95.840 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 89.120 4.000 89.720 ;
=======
        RECT 0.000 100.680 4.000 101.280 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 93.880 4.000 94.480 ;
=======
        RECT 0.000 106.120 4.000 106.720 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 6.840 4.000 7.440 ;
=======
        RECT 0.000 8.200 4.000 8.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 98.640 4.000 99.240 ;
=======
        RECT 0.000 111.560 4.000 112.160 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 103.400 4.000 104.000 ;
=======
        RECT 0.000 117.000 4.000 117.600 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 108.160 4.000 108.760 ;
=======
        RECT 0.000 122.440 4.000 123.040 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 112.920 4.000 113.520 ;
=======
        RECT 0.000 127.880 4.000 128.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 117.680 4.000 118.280 ;
=======
        RECT 0.000 133.320 4.000 133.920 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 122.440 4.000 123.040 ;
=======
        RECT 0.000 138.760 4.000 139.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 127.200 4.000 127.800 ;
=======
        RECT 0.000 144.200 4.000 144.800 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 132.640 4.000 133.240 ;
=======
        RECT 0.000 149.640 4.000 150.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 137.400 4.000 138.000 ;
=======
        RECT 0.000 155.080 4.000 155.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 142.160 4.000 142.760 ;
=======
        RECT 0.000 160.520 4.000 161.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 11.600 4.000 12.200 ;
=======
        RECT 0.000 13.640 4.000 14.240 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 146.920 4.000 147.520 ;
=======
        RECT 0.000 165.960 4.000 166.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 151.680 4.000 152.280 ;
=======
        RECT 0.000 171.400 4.000 172.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 16.360 4.000 16.960 ;
=======
        RECT 0.000 19.080 4.000 19.680 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 21.120 4.000 21.720 ;
=======
        RECT 0.000 24.520 4.000 25.120 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 25.880 4.000 26.480 ;
=======
        RECT 0.000 29.960 4.000 30.560 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 30.640 4.000 31.240 ;
=======
        RECT 0.000 35.400 4.000 36.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 35.400 4.000 36.000 ;
=======
        RECT 0.000 40.840 4.000 41.440 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 40.160 4.000 40.760 ;
=======
        RECT 0.000 46.280 4.000 46.880 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
<<<<<<< HEAD
        RECT 0.000 45.600 4.000 46.200 ;
=======
        RECT 0.000 51.720 4.000 52.320 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 23.550 296.000 23.830 300.000 ;
=======
        RECT 22.170 296.000 22.450 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 26.310 296.000 26.590 300.000 ;
=======
        RECT 25.390 296.000 25.670 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 29.530 296.000 29.810 300.000 ;
=======
        RECT 28.150 296.000 28.430 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 32.750 296.000 33.030 300.000 ;
=======
        RECT 31.370 296.000 31.650 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 296.000 7.730 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
<<<<<<< HEAD
        RECT 13.890 296.000 14.170 300.000 ;
=======
        RECT 13.430 296.000 13.710 300.000 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
<<<<<<< HEAD
        RECT 5.520 10.795 296.095 288.405 ;
      LAYER met1 ;
        RECT 1.450 6.500 296.155 289.300 ;
      LAYER met2 ;
        RECT 2.030 295.720 3.950 298.365 ;
        RECT 4.790 295.720 7.170 298.365 ;
        RECT 8.010 295.720 10.390 298.365 ;
        RECT 11.230 295.720 13.610 298.365 ;
        RECT 14.450 295.720 16.830 298.365 ;
        RECT 17.670 295.720 20.050 298.365 ;
        RECT 20.890 295.720 23.270 298.365 ;
        RECT 24.110 295.720 26.030 298.365 ;
        RECT 26.870 295.720 29.250 298.365 ;
        RECT 30.090 295.720 32.470 298.365 ;
        RECT 33.310 295.720 35.690 298.365 ;
        RECT 36.530 295.720 38.910 298.365 ;
        RECT 39.750 295.720 42.130 298.365 ;
        RECT 42.970 295.720 45.350 298.365 ;
        RECT 46.190 295.720 48.110 298.365 ;
        RECT 48.950 295.720 51.330 298.365 ;
        RECT 52.170 295.720 54.550 298.365 ;
        RECT 55.390 295.720 57.770 298.365 ;
        RECT 58.610 295.720 60.990 298.365 ;
        RECT 61.830 295.720 64.210 298.365 ;
        RECT 65.050 295.720 67.430 298.365 ;
        RECT 68.270 295.720 70.190 298.365 ;
        RECT 71.030 295.720 73.410 298.365 ;
        RECT 74.250 295.720 76.630 298.365 ;
        RECT 77.470 295.720 79.850 298.365 ;
        RECT 80.690 295.720 83.070 298.365 ;
        RECT 83.910 295.720 86.290 298.365 ;
        RECT 87.130 295.720 89.510 298.365 ;
        RECT 90.350 295.720 92.730 298.365 ;
        RECT 93.570 295.720 95.490 298.365 ;
        RECT 96.330 295.720 98.710 298.365 ;
        RECT 99.550 295.720 101.930 298.365 ;
        RECT 102.770 295.720 105.150 298.365 ;
        RECT 105.990 295.720 108.370 298.365 ;
        RECT 109.210 295.720 111.590 298.365 ;
        RECT 112.430 295.720 114.810 298.365 ;
        RECT 115.650 295.720 117.570 298.365 ;
        RECT 118.410 295.720 120.790 298.365 ;
        RECT 121.630 295.720 124.010 298.365 ;
        RECT 124.850 295.720 127.230 298.365 ;
        RECT 128.070 295.720 130.450 298.365 ;
        RECT 131.290 295.720 133.670 298.365 ;
        RECT 134.510 295.720 136.890 298.365 ;
        RECT 137.730 295.720 139.650 298.365 ;
        RECT 140.490 295.720 142.870 298.365 ;
        RECT 143.710 295.720 146.090 298.365 ;
        RECT 146.930 295.720 149.310 298.365 ;
        RECT 150.150 295.720 152.530 298.365 ;
        RECT 153.370 295.720 155.750 298.365 ;
        RECT 156.590 295.720 158.970 298.365 ;
        RECT 159.810 295.720 162.190 298.365 ;
        RECT 163.030 295.720 164.950 298.365 ;
        RECT 165.790 295.720 168.170 298.365 ;
        RECT 169.010 295.720 171.390 298.365 ;
        RECT 172.230 295.720 174.610 298.365 ;
        RECT 175.450 295.720 177.830 298.365 ;
        RECT 178.670 295.720 181.050 298.365 ;
        RECT 181.890 295.720 184.270 298.365 ;
        RECT 185.110 295.720 187.030 298.365 ;
        RECT 187.870 295.720 190.250 298.365 ;
        RECT 191.090 295.720 193.470 298.365 ;
        RECT 194.310 295.720 196.690 298.365 ;
        RECT 197.530 295.720 199.910 298.365 ;
        RECT 200.750 295.720 203.130 298.365 ;
        RECT 203.970 295.720 206.350 298.365 ;
        RECT 207.190 295.720 209.110 298.365 ;
        RECT 209.950 295.720 212.330 298.365 ;
        RECT 213.170 295.720 215.550 298.365 ;
        RECT 216.390 295.720 218.770 298.365 ;
        RECT 219.610 295.720 221.990 298.365 ;
        RECT 222.830 295.720 225.210 298.365 ;
        RECT 226.050 295.720 228.430 298.365 ;
        RECT 229.270 295.720 231.650 298.365 ;
        RECT 232.490 295.720 234.410 298.365 ;
        RECT 235.250 295.720 237.630 298.365 ;
        RECT 238.470 295.720 240.850 298.365 ;
        RECT 241.690 295.720 244.070 298.365 ;
        RECT 244.910 295.720 247.290 298.365 ;
        RECT 248.130 295.720 250.510 298.365 ;
        RECT 251.350 295.720 253.730 298.365 ;
        RECT 254.570 295.720 256.490 298.365 ;
        RECT 257.330 295.720 259.710 298.365 ;
        RECT 260.550 295.720 262.930 298.365 ;
        RECT 263.770 295.720 266.150 298.365 ;
        RECT 266.990 295.720 269.370 298.365 ;
        RECT 270.210 295.720 272.590 298.365 ;
        RECT 273.430 295.720 275.810 298.365 ;
        RECT 276.650 295.720 278.570 298.365 ;
        RECT 279.410 295.720 281.790 298.365 ;
        RECT 282.630 295.720 285.010 298.365 ;
        RECT 285.850 295.720 288.230 298.365 ;
        RECT 289.070 295.720 291.450 298.365 ;
        RECT 292.290 295.720 294.670 298.365 ;
        RECT 1.480 4.280 295.220 295.720 ;
        RECT 1.480 0.270 8.090 4.280 ;
        RECT 8.930 0.270 24.650 4.280 ;
        RECT 25.490 0.270 41.210 4.280 ;
        RECT 42.050 0.270 57.770 4.280 ;
        RECT 58.610 0.270 74.330 4.280 ;
        RECT 75.170 0.270 91.350 4.280 ;
        RECT 92.190 0.270 107.910 4.280 ;
        RECT 108.750 0.270 124.470 4.280 ;
        RECT 125.310 0.270 141.030 4.280 ;
        RECT 141.870 0.270 158.050 4.280 ;
        RECT 158.890 0.270 174.610 4.280 ;
        RECT 175.450 0.270 191.170 4.280 ;
        RECT 192.010 0.270 207.730 4.280 ;
        RECT 208.570 0.270 224.290 4.280 ;
        RECT 225.130 0.270 241.310 4.280 ;
        RECT 242.150 0.270 257.870 4.280 ;
        RECT 258.710 0.270 274.430 4.280 ;
        RECT 275.270 0.270 290.990 4.280 ;
        RECT 291.830 0.270 295.220 4.280 ;
      LAYER met3 ;
        RECT 4.000 297.520 295.600 298.345 ;
        RECT 4.400 297.480 295.600 297.520 ;
        RECT 4.400 296.840 296.000 297.480 ;
        RECT 4.400 296.120 295.600 296.840 ;
        RECT 4.000 295.440 295.600 296.120 ;
        RECT 4.000 294.800 296.000 295.440 ;
        RECT 4.000 293.400 295.600 294.800 ;
        RECT 4.000 292.760 296.000 293.400 ;
        RECT 4.400 291.360 295.600 292.760 ;
        RECT 4.000 290.720 296.000 291.360 ;
        RECT 4.000 289.320 295.600 290.720 ;
        RECT 4.000 288.680 296.000 289.320 ;
        RECT 4.000 288.000 295.600 288.680 ;
        RECT 4.400 287.280 295.600 288.000 ;
        RECT 4.400 286.640 296.000 287.280 ;
        RECT 4.400 286.600 295.600 286.640 ;
        RECT 4.000 285.240 295.600 286.600 ;
        RECT 4.000 284.600 296.000 285.240 ;
        RECT 4.000 283.240 295.600 284.600 ;
        RECT 4.400 283.200 295.600 283.240 ;
        RECT 4.400 282.560 296.000 283.200 ;
        RECT 4.400 281.840 295.600 282.560 ;
        RECT 4.000 281.160 295.600 281.840 ;
        RECT 4.000 280.520 296.000 281.160 ;
        RECT 4.000 279.120 295.600 280.520 ;
        RECT 4.000 278.480 296.000 279.120 ;
        RECT 4.400 277.080 295.600 278.480 ;
        RECT 4.000 276.440 296.000 277.080 ;
        RECT 4.000 275.040 295.600 276.440 ;
        RECT 4.000 274.400 296.000 275.040 ;
        RECT 4.000 273.720 295.600 274.400 ;
        RECT 4.400 273.000 295.600 273.720 ;
        RECT 4.400 272.360 296.000 273.000 ;
        RECT 4.400 272.320 295.600 272.360 ;
        RECT 4.000 270.960 295.600 272.320 ;
        RECT 4.000 270.320 296.000 270.960 ;
        RECT 4.000 268.960 295.600 270.320 ;
        RECT 4.400 268.920 295.600 268.960 ;
        RECT 4.400 268.280 296.000 268.920 ;
        RECT 4.400 267.560 295.600 268.280 ;
        RECT 4.000 266.880 295.600 267.560 ;
        RECT 4.000 266.240 296.000 266.880 ;
        RECT 4.000 264.840 295.600 266.240 ;
        RECT 4.000 264.200 296.000 264.840 ;
        RECT 4.400 262.800 295.600 264.200 ;
        RECT 4.000 262.160 296.000 262.800 ;
        RECT 4.000 260.760 295.600 262.160 ;
        RECT 4.000 260.120 296.000 260.760 ;
        RECT 4.000 258.760 295.600 260.120 ;
        RECT 4.400 258.720 295.600 258.760 ;
        RECT 4.400 258.080 296.000 258.720 ;
        RECT 4.400 257.360 295.600 258.080 ;
        RECT 4.000 256.680 295.600 257.360 ;
        RECT 4.000 256.040 296.000 256.680 ;
=======
        RECT 5.520 10.795 296.555 288.405 ;
      LAYER met1 ;
        RECT 1.450 10.240 296.615 289.640 ;
      LAYER met2 ;
        RECT 2.030 295.720 3.950 296.210 ;
        RECT 4.790 295.720 7.170 296.210 ;
        RECT 8.010 295.720 9.930 296.210 ;
        RECT 10.770 295.720 13.150 296.210 ;
        RECT 13.990 295.720 15.910 296.210 ;
        RECT 16.750 295.720 19.130 296.210 ;
        RECT 19.970 295.720 21.890 296.210 ;
        RECT 22.730 295.720 25.110 296.210 ;
        RECT 25.950 295.720 27.870 296.210 ;
        RECT 28.710 295.720 31.090 296.210 ;
        RECT 31.930 295.720 33.850 296.210 ;
        RECT 34.690 295.720 37.070 296.210 ;
        RECT 37.910 295.720 39.830 296.210 ;
        RECT 40.670 295.720 43.050 296.210 ;
        RECT 43.890 295.720 45.810 296.210 ;
        RECT 46.650 295.720 49.030 296.210 ;
        RECT 49.870 295.720 51.790 296.210 ;
        RECT 52.630 295.720 55.010 296.210 ;
        RECT 55.850 295.720 57.770 296.210 ;
        RECT 58.610 295.720 60.990 296.210 ;
        RECT 61.830 295.720 63.750 296.210 ;
        RECT 64.590 295.720 66.970 296.210 ;
        RECT 67.810 295.720 69.730 296.210 ;
        RECT 70.570 295.720 72.950 296.210 ;
        RECT 73.790 295.720 76.170 296.210 ;
        RECT 77.010 295.720 78.930 296.210 ;
        RECT 79.770 295.720 82.150 296.210 ;
        RECT 82.990 295.720 84.910 296.210 ;
        RECT 85.750 295.720 88.130 296.210 ;
        RECT 88.970 295.720 90.890 296.210 ;
        RECT 91.730 295.720 94.110 296.210 ;
        RECT 94.950 295.720 96.870 296.210 ;
        RECT 97.710 295.720 100.090 296.210 ;
        RECT 100.930 295.720 102.850 296.210 ;
        RECT 103.690 295.720 106.070 296.210 ;
        RECT 106.910 295.720 108.830 296.210 ;
        RECT 109.670 295.720 112.050 296.210 ;
        RECT 112.890 295.720 114.810 296.210 ;
        RECT 115.650 295.720 118.030 296.210 ;
        RECT 118.870 295.720 120.790 296.210 ;
        RECT 121.630 295.720 124.010 296.210 ;
        RECT 124.850 295.720 126.770 296.210 ;
        RECT 127.610 295.720 129.990 296.210 ;
        RECT 130.830 295.720 132.750 296.210 ;
        RECT 133.590 295.720 135.970 296.210 ;
        RECT 136.810 295.720 138.730 296.210 ;
        RECT 139.570 295.720 141.950 296.210 ;
        RECT 142.790 295.720 144.710 296.210 ;
        RECT 145.550 295.720 147.930 296.210 ;
        RECT 148.770 295.720 151.150 296.210 ;
        RECT 151.990 295.720 153.910 296.210 ;
        RECT 154.750 295.720 157.130 296.210 ;
        RECT 157.970 295.720 159.890 296.210 ;
        RECT 160.730 295.720 163.110 296.210 ;
        RECT 163.950 295.720 165.870 296.210 ;
        RECT 166.710 295.720 169.090 296.210 ;
        RECT 169.930 295.720 171.850 296.210 ;
        RECT 172.690 295.720 175.070 296.210 ;
        RECT 175.910 295.720 177.830 296.210 ;
        RECT 178.670 295.720 181.050 296.210 ;
        RECT 181.890 295.720 183.810 296.210 ;
        RECT 184.650 295.720 187.030 296.210 ;
        RECT 187.870 295.720 189.790 296.210 ;
        RECT 190.630 295.720 193.010 296.210 ;
        RECT 193.850 295.720 195.770 296.210 ;
        RECT 196.610 295.720 198.990 296.210 ;
        RECT 199.830 295.720 201.750 296.210 ;
        RECT 202.590 295.720 204.970 296.210 ;
        RECT 205.810 295.720 207.730 296.210 ;
        RECT 208.570 295.720 210.950 296.210 ;
        RECT 211.790 295.720 213.710 296.210 ;
        RECT 214.550 295.720 216.930 296.210 ;
        RECT 217.770 295.720 219.690 296.210 ;
        RECT 220.530 295.720 222.910 296.210 ;
        RECT 223.750 295.720 226.130 296.210 ;
        RECT 226.970 295.720 228.890 296.210 ;
        RECT 229.730 295.720 232.110 296.210 ;
        RECT 232.950 295.720 234.870 296.210 ;
        RECT 235.710 295.720 238.090 296.210 ;
        RECT 238.930 295.720 240.850 296.210 ;
        RECT 241.690 295.720 244.070 296.210 ;
        RECT 244.910 295.720 246.830 296.210 ;
        RECT 247.670 295.720 250.050 296.210 ;
        RECT 250.890 295.720 252.810 296.210 ;
        RECT 253.650 295.720 256.030 296.210 ;
        RECT 256.870 295.720 258.790 296.210 ;
        RECT 259.630 295.720 262.010 296.210 ;
        RECT 262.850 295.720 264.770 296.210 ;
        RECT 265.610 295.720 267.990 296.210 ;
        RECT 268.830 295.720 270.750 296.210 ;
        RECT 271.590 295.720 273.970 296.210 ;
        RECT 274.810 295.720 276.730 296.210 ;
        RECT 277.570 295.720 279.950 296.210 ;
        RECT 280.790 295.720 282.710 296.210 ;
        RECT 283.550 295.720 285.930 296.210 ;
        RECT 286.770 295.720 288.690 296.210 ;
        RECT 289.530 295.720 291.910 296.210 ;
        RECT 292.750 295.720 293.840 296.210 ;
        RECT 1.480 4.280 293.840 295.720 ;
        RECT 1.480 2.875 5.790 4.280 ;
        RECT 6.630 2.875 17.750 4.280 ;
        RECT 18.590 2.875 29.710 4.280 ;
        RECT 30.550 2.875 41.670 4.280 ;
        RECT 42.510 2.875 53.630 4.280 ;
        RECT 54.470 2.875 65.590 4.280 ;
        RECT 66.430 2.875 77.550 4.280 ;
        RECT 78.390 2.875 89.510 4.280 ;
        RECT 90.350 2.875 101.470 4.280 ;
        RECT 102.310 2.875 113.430 4.280 ;
        RECT 114.270 2.875 125.390 4.280 ;
        RECT 126.230 2.875 137.350 4.280 ;
        RECT 138.190 2.875 149.310 4.280 ;
        RECT 150.150 2.875 161.730 4.280 ;
        RECT 162.570 2.875 173.690 4.280 ;
        RECT 174.530 2.875 185.650 4.280 ;
        RECT 186.490 2.875 197.610 4.280 ;
        RECT 198.450 2.875 209.570 4.280 ;
        RECT 210.410 2.875 221.530 4.280 ;
        RECT 222.370 2.875 233.490 4.280 ;
        RECT 234.330 2.875 245.450 4.280 ;
        RECT 246.290 2.875 257.410 4.280 ;
        RECT 258.250 2.875 269.370 4.280 ;
        RECT 270.210 2.875 281.330 4.280 ;
        RECT 282.170 2.875 293.290 4.280 ;
      LAYER met3 ;
        RECT 4.400 291.360 295.600 291.545 ;
        RECT 4.400 290.720 296.000 291.360 ;
        RECT 4.400 290.680 295.600 290.720 ;
        RECT 4.000 289.320 295.600 290.680 ;
        RECT 4.000 288.680 296.000 289.320 ;
        RECT 4.000 287.280 295.600 288.680 ;
        RECT 4.000 286.640 296.000 287.280 ;
        RECT 4.400 285.960 296.000 286.640 ;
        RECT 4.400 285.240 295.600 285.960 ;
        RECT 4.000 284.560 295.600 285.240 ;
        RECT 4.000 283.920 296.000 284.560 ;
        RECT 4.000 282.520 295.600 283.920 ;
        RECT 4.000 281.880 296.000 282.520 ;
        RECT 4.000 281.200 295.600 281.880 ;
        RECT 4.400 280.480 295.600 281.200 ;
        RECT 4.400 279.840 296.000 280.480 ;
        RECT 4.400 279.800 295.600 279.840 ;
        RECT 4.000 278.440 295.600 279.800 ;
        RECT 4.000 277.800 296.000 278.440 ;
        RECT 4.000 276.400 295.600 277.800 ;
        RECT 4.000 275.760 296.000 276.400 ;
        RECT 4.400 274.360 295.600 275.760 ;
        RECT 4.000 273.720 296.000 274.360 ;
        RECT 4.000 272.320 295.600 273.720 ;
        RECT 4.000 271.000 296.000 272.320 ;
        RECT 4.000 270.320 295.600 271.000 ;
        RECT 4.400 269.600 295.600 270.320 ;
        RECT 4.400 268.960 296.000 269.600 ;
        RECT 4.400 268.920 295.600 268.960 ;
        RECT 4.000 267.560 295.600 268.920 ;
        RECT 4.000 266.920 296.000 267.560 ;
        RECT 4.000 265.520 295.600 266.920 ;
        RECT 4.000 264.880 296.000 265.520 ;
        RECT 4.400 263.480 295.600 264.880 ;
        RECT 4.000 262.840 296.000 263.480 ;
        RECT 4.000 261.440 295.600 262.840 ;
        RECT 4.000 260.800 296.000 261.440 ;
        RECT 4.000 259.440 295.600 260.800 ;
        RECT 4.400 259.400 295.600 259.440 ;
        RECT 4.400 258.760 296.000 259.400 ;
        RECT 4.400 258.040 295.600 258.760 ;
        RECT 4.000 257.360 295.600 258.040 ;
        RECT 4.000 256.040 296.000 257.360 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
        RECT 4.000 254.640 295.600 256.040 ;
        RECT 4.000 254.000 296.000 254.640 ;
        RECT 4.400 252.600 295.600 254.000 ;
        RECT 4.000 251.960 296.000 252.600 ;
        RECT 4.000 250.560 295.600 251.960 ;
<<<<<<< HEAD
        RECT 4.000 249.240 296.000 250.560 ;
        RECT 4.400 247.840 295.600 249.240 ;
        RECT 4.000 247.200 296.000 247.840 ;
        RECT 4.000 245.800 295.600 247.200 ;
        RECT 4.000 245.160 296.000 245.800 ;
        RECT 4.000 244.480 295.600 245.160 ;
        RECT 4.400 243.760 295.600 244.480 ;
        RECT 4.400 243.120 296.000 243.760 ;
        RECT 4.400 243.080 295.600 243.120 ;
        RECT 4.000 241.720 295.600 243.080 ;
        RECT 4.000 241.080 296.000 241.720 ;
        RECT 4.000 239.720 295.600 241.080 ;
        RECT 4.400 239.680 295.600 239.720 ;
        RECT 4.400 239.040 296.000 239.680 ;
        RECT 4.400 238.320 295.600 239.040 ;
        RECT 4.000 237.640 295.600 238.320 ;
        RECT 4.000 237.000 296.000 237.640 ;
        RECT 4.000 235.600 295.600 237.000 ;
        RECT 4.000 234.960 296.000 235.600 ;
        RECT 4.400 233.560 295.600 234.960 ;
        RECT 4.000 232.920 296.000 233.560 ;
        RECT 4.000 231.520 295.600 232.920 ;
        RECT 4.000 230.880 296.000 231.520 ;
        RECT 4.000 230.200 295.600 230.880 ;
        RECT 4.400 229.480 295.600 230.200 ;
        RECT 4.400 228.840 296.000 229.480 ;
        RECT 4.400 228.800 295.600 228.840 ;
        RECT 4.000 227.440 295.600 228.800 ;
        RECT 4.000 226.800 296.000 227.440 ;
        RECT 4.000 225.440 295.600 226.800 ;
        RECT 4.400 225.400 295.600 225.440 ;
        RECT 4.400 224.760 296.000 225.400 ;
        RECT 4.400 224.040 295.600 224.760 ;
        RECT 4.000 223.360 295.600 224.040 ;
        RECT 4.000 222.720 296.000 223.360 ;
        RECT 4.000 221.320 295.600 222.720 ;
        RECT 4.000 220.680 296.000 221.320 ;
        RECT 4.400 219.280 295.600 220.680 ;
        RECT 4.000 218.640 296.000 219.280 ;
        RECT 4.000 217.240 295.600 218.640 ;
        RECT 4.000 216.600 296.000 217.240 ;
        RECT 4.000 215.240 295.600 216.600 ;
        RECT 4.400 215.200 295.600 215.240 ;
        RECT 4.400 214.560 296.000 215.200 ;
        RECT 4.400 213.840 295.600 214.560 ;
        RECT 4.000 213.160 295.600 213.840 ;
        RECT 4.000 212.520 296.000 213.160 ;
        RECT 4.000 211.120 295.600 212.520 ;
        RECT 4.000 210.480 296.000 211.120 ;
        RECT 4.400 209.080 295.600 210.480 ;
        RECT 4.000 208.440 296.000 209.080 ;
        RECT 4.000 207.040 295.600 208.440 ;
        RECT 4.000 206.400 296.000 207.040 ;
        RECT 4.000 205.720 295.600 206.400 ;
        RECT 4.400 205.000 295.600 205.720 ;
        RECT 4.400 204.360 296.000 205.000 ;
        RECT 4.400 204.320 295.600 204.360 ;
        RECT 4.000 202.960 295.600 204.320 ;
        RECT 4.000 202.320 296.000 202.960 ;
        RECT 4.000 200.960 295.600 202.320 ;
        RECT 4.400 200.920 295.600 200.960 ;
        RECT 4.400 199.600 296.000 200.920 ;
        RECT 4.400 199.560 295.600 199.600 ;
        RECT 4.000 198.200 295.600 199.560 ;
        RECT 4.000 197.560 296.000 198.200 ;
        RECT 4.000 196.200 295.600 197.560 ;
        RECT 4.400 196.160 295.600 196.200 ;
        RECT 4.400 195.520 296.000 196.160 ;
        RECT 4.400 194.800 295.600 195.520 ;
        RECT 4.000 194.120 295.600 194.800 ;
        RECT 4.000 193.480 296.000 194.120 ;
        RECT 4.000 192.080 295.600 193.480 ;
        RECT 4.000 191.440 296.000 192.080 ;
        RECT 4.400 190.040 295.600 191.440 ;
        RECT 4.000 189.400 296.000 190.040 ;
        RECT 4.000 188.000 295.600 189.400 ;
        RECT 4.000 187.360 296.000 188.000 ;
        RECT 4.000 186.680 295.600 187.360 ;
        RECT 4.400 185.960 295.600 186.680 ;
        RECT 4.400 185.320 296.000 185.960 ;
        RECT 4.400 185.280 295.600 185.320 ;
        RECT 4.000 183.920 295.600 185.280 ;
        RECT 4.000 183.280 296.000 183.920 ;
        RECT 4.000 181.920 295.600 183.280 ;
        RECT 4.400 181.880 295.600 181.920 ;
        RECT 4.400 181.240 296.000 181.880 ;
        RECT 4.400 180.520 295.600 181.240 ;
        RECT 4.000 179.840 295.600 180.520 ;
        RECT 4.000 179.200 296.000 179.840 ;
        RECT 4.000 177.800 295.600 179.200 ;
        RECT 4.000 177.160 296.000 177.800 ;
        RECT 4.400 175.760 295.600 177.160 ;
        RECT 4.000 175.120 296.000 175.760 ;
        RECT 4.000 173.720 295.600 175.120 ;
        RECT 4.000 173.080 296.000 173.720 ;
        RECT 4.000 171.720 295.600 173.080 ;
        RECT 4.400 171.680 295.600 171.720 ;
        RECT 4.400 171.040 296.000 171.680 ;
        RECT 4.400 170.320 295.600 171.040 ;
        RECT 4.000 169.640 295.600 170.320 ;
        RECT 4.000 169.000 296.000 169.640 ;
        RECT 4.000 167.600 295.600 169.000 ;
        RECT 4.000 166.960 296.000 167.600 ;
        RECT 4.400 165.560 295.600 166.960 ;
        RECT 4.000 164.920 296.000 165.560 ;
        RECT 4.000 163.520 295.600 164.920 ;
        RECT 4.000 162.880 296.000 163.520 ;
        RECT 4.000 162.200 295.600 162.880 ;
        RECT 4.400 161.480 295.600 162.200 ;
        RECT 4.400 160.840 296.000 161.480 ;
        RECT 4.400 160.800 295.600 160.840 ;
        RECT 4.000 159.440 295.600 160.800 ;
        RECT 4.000 158.800 296.000 159.440 ;
        RECT 4.000 157.440 295.600 158.800 ;
        RECT 4.400 157.400 295.600 157.440 ;
        RECT 4.400 156.760 296.000 157.400 ;
        RECT 4.400 156.040 295.600 156.760 ;
        RECT 4.000 155.360 295.600 156.040 ;
        RECT 4.000 154.720 296.000 155.360 ;
        RECT 4.000 153.320 295.600 154.720 ;
        RECT 4.000 152.680 296.000 153.320 ;
        RECT 4.400 151.280 295.600 152.680 ;
        RECT 4.000 149.960 296.000 151.280 ;
        RECT 4.000 148.560 295.600 149.960 ;
        RECT 4.000 147.920 296.000 148.560 ;
        RECT 4.400 146.520 295.600 147.920 ;
        RECT 4.000 145.880 296.000 146.520 ;
        RECT 4.000 144.480 295.600 145.880 ;
        RECT 4.000 143.840 296.000 144.480 ;
        RECT 4.000 143.160 295.600 143.840 ;
        RECT 4.400 142.440 295.600 143.160 ;
        RECT 4.400 141.800 296.000 142.440 ;
        RECT 4.400 141.760 295.600 141.800 ;
        RECT 4.000 140.400 295.600 141.760 ;
        RECT 4.000 139.760 296.000 140.400 ;
        RECT 4.000 138.400 295.600 139.760 ;
        RECT 4.400 138.360 295.600 138.400 ;
        RECT 4.400 137.720 296.000 138.360 ;
        RECT 4.400 137.000 295.600 137.720 ;
        RECT 4.000 136.320 295.600 137.000 ;
        RECT 4.000 135.680 296.000 136.320 ;
        RECT 4.000 134.280 295.600 135.680 ;
        RECT 4.000 133.640 296.000 134.280 ;
        RECT 4.400 132.240 295.600 133.640 ;
        RECT 4.000 131.600 296.000 132.240 ;
        RECT 4.000 130.200 295.600 131.600 ;
        RECT 4.000 129.560 296.000 130.200 ;
        RECT 4.000 128.200 295.600 129.560 ;
        RECT 4.400 128.160 295.600 128.200 ;
        RECT 4.400 127.520 296.000 128.160 ;
        RECT 4.400 126.800 295.600 127.520 ;
        RECT 4.000 126.120 295.600 126.800 ;
=======
        RECT 4.000 249.920 296.000 250.560 ;
        RECT 4.000 248.560 295.600 249.920 ;
        RECT 4.400 248.520 295.600 248.560 ;
        RECT 4.400 247.880 296.000 248.520 ;
        RECT 4.400 247.160 295.600 247.880 ;
        RECT 4.000 246.480 295.600 247.160 ;
        RECT 4.000 245.840 296.000 246.480 ;
        RECT 4.000 244.440 295.600 245.840 ;
        RECT 4.000 243.120 296.000 244.440 ;
        RECT 4.400 241.720 295.600 243.120 ;
        RECT 4.000 241.080 296.000 241.720 ;
        RECT 4.000 239.680 295.600 241.080 ;
        RECT 4.000 239.040 296.000 239.680 ;
        RECT 4.000 237.680 295.600 239.040 ;
        RECT 4.400 237.640 295.600 237.680 ;
        RECT 4.400 237.000 296.000 237.640 ;
        RECT 4.400 236.280 295.600 237.000 ;
        RECT 4.000 235.600 295.600 236.280 ;
        RECT 4.000 234.960 296.000 235.600 ;
        RECT 4.000 233.560 295.600 234.960 ;
        RECT 4.000 232.920 296.000 233.560 ;
        RECT 4.000 232.240 295.600 232.920 ;
        RECT 4.400 231.520 295.600 232.240 ;
        RECT 4.400 230.880 296.000 231.520 ;
        RECT 4.400 230.840 295.600 230.880 ;
        RECT 4.000 229.480 295.600 230.840 ;
        RECT 4.000 228.160 296.000 229.480 ;
        RECT 4.000 226.800 295.600 228.160 ;
        RECT 4.400 226.760 295.600 226.800 ;
        RECT 4.400 226.120 296.000 226.760 ;
        RECT 4.400 225.400 295.600 226.120 ;
        RECT 4.000 224.720 295.600 225.400 ;
        RECT 4.000 224.080 296.000 224.720 ;
        RECT 4.000 222.680 295.600 224.080 ;
        RECT 4.000 222.040 296.000 222.680 ;
        RECT 4.000 221.360 295.600 222.040 ;
        RECT 4.400 220.640 295.600 221.360 ;
        RECT 4.400 220.000 296.000 220.640 ;
        RECT 4.400 219.960 295.600 220.000 ;
        RECT 4.000 218.600 295.600 219.960 ;
        RECT 4.000 217.960 296.000 218.600 ;
        RECT 4.000 216.560 295.600 217.960 ;
        RECT 4.000 215.920 296.000 216.560 ;
        RECT 4.400 214.520 295.600 215.920 ;
        RECT 4.000 213.200 296.000 214.520 ;
        RECT 4.000 211.800 295.600 213.200 ;
        RECT 4.000 211.160 296.000 211.800 ;
        RECT 4.000 210.480 295.600 211.160 ;
        RECT 4.400 209.760 295.600 210.480 ;
        RECT 4.400 209.120 296.000 209.760 ;
        RECT 4.400 209.080 295.600 209.120 ;
        RECT 4.000 207.720 295.600 209.080 ;
        RECT 4.000 207.080 296.000 207.720 ;
        RECT 4.000 205.680 295.600 207.080 ;
        RECT 4.000 205.040 296.000 205.680 ;
        RECT 4.400 203.640 295.600 205.040 ;
        RECT 4.000 203.000 296.000 203.640 ;
        RECT 4.000 201.600 295.600 203.000 ;
        RECT 4.000 200.280 296.000 201.600 ;
        RECT 4.000 199.600 295.600 200.280 ;
        RECT 4.400 198.880 295.600 199.600 ;
        RECT 4.400 198.240 296.000 198.880 ;
        RECT 4.400 198.200 295.600 198.240 ;
        RECT 4.000 196.840 295.600 198.200 ;
        RECT 4.000 196.200 296.000 196.840 ;
        RECT 4.000 194.800 295.600 196.200 ;
        RECT 4.000 194.160 296.000 194.800 ;
        RECT 4.400 192.760 295.600 194.160 ;
        RECT 4.000 192.120 296.000 192.760 ;
        RECT 4.000 190.720 295.600 192.120 ;
        RECT 4.000 190.080 296.000 190.720 ;
        RECT 4.000 188.720 295.600 190.080 ;
        RECT 4.400 188.680 295.600 188.720 ;
        RECT 4.400 188.040 296.000 188.680 ;
        RECT 4.400 187.320 295.600 188.040 ;
        RECT 4.000 186.640 295.600 187.320 ;
        RECT 4.000 185.320 296.000 186.640 ;
        RECT 4.000 183.920 295.600 185.320 ;
        RECT 4.000 183.280 296.000 183.920 ;
        RECT 4.400 181.880 295.600 183.280 ;
        RECT 4.000 181.240 296.000 181.880 ;
        RECT 4.000 179.840 295.600 181.240 ;
        RECT 4.000 179.200 296.000 179.840 ;
        RECT 4.000 177.840 295.600 179.200 ;
        RECT 4.400 177.800 295.600 177.840 ;
        RECT 4.400 177.160 296.000 177.800 ;
        RECT 4.400 176.440 295.600 177.160 ;
        RECT 4.000 175.760 295.600 176.440 ;
        RECT 4.000 175.120 296.000 175.760 ;
        RECT 4.000 173.720 295.600 175.120 ;
        RECT 4.000 173.080 296.000 173.720 ;
        RECT 4.000 172.400 295.600 173.080 ;
        RECT 4.400 171.680 295.600 172.400 ;
        RECT 4.400 171.000 296.000 171.680 ;
        RECT 4.000 170.360 296.000 171.000 ;
        RECT 4.000 168.960 295.600 170.360 ;
        RECT 4.000 168.320 296.000 168.960 ;
        RECT 4.000 166.960 295.600 168.320 ;
        RECT 4.400 166.920 295.600 166.960 ;
        RECT 4.400 166.280 296.000 166.920 ;
        RECT 4.400 165.560 295.600 166.280 ;
        RECT 4.000 164.880 295.600 165.560 ;
        RECT 4.000 164.240 296.000 164.880 ;
        RECT 4.000 162.840 295.600 164.240 ;
        RECT 4.000 162.200 296.000 162.840 ;
        RECT 4.000 161.520 295.600 162.200 ;
        RECT 4.400 160.800 295.600 161.520 ;
        RECT 4.400 160.160 296.000 160.800 ;
        RECT 4.400 160.120 295.600 160.160 ;
        RECT 4.000 158.760 295.600 160.120 ;
        RECT 4.000 157.440 296.000 158.760 ;
        RECT 4.000 156.080 295.600 157.440 ;
        RECT 4.400 156.040 295.600 156.080 ;
        RECT 4.400 155.400 296.000 156.040 ;
        RECT 4.400 154.680 295.600 155.400 ;
        RECT 4.000 154.000 295.600 154.680 ;
        RECT 4.000 153.360 296.000 154.000 ;
        RECT 4.000 151.960 295.600 153.360 ;
        RECT 4.000 151.320 296.000 151.960 ;
        RECT 4.000 150.640 295.600 151.320 ;
        RECT 4.400 149.920 295.600 150.640 ;
        RECT 4.400 149.280 296.000 149.920 ;
        RECT 4.400 149.240 295.600 149.280 ;
        RECT 4.000 147.880 295.600 149.240 ;
        RECT 4.000 147.240 296.000 147.880 ;
        RECT 4.000 145.840 295.600 147.240 ;
        RECT 4.000 145.200 296.000 145.840 ;
        RECT 4.400 143.800 295.600 145.200 ;
        RECT 4.000 142.480 296.000 143.800 ;
        RECT 4.000 141.080 295.600 142.480 ;
        RECT 4.000 140.440 296.000 141.080 ;
        RECT 4.000 139.760 295.600 140.440 ;
        RECT 4.400 139.040 295.600 139.760 ;
        RECT 4.400 138.400 296.000 139.040 ;
        RECT 4.400 138.360 295.600 138.400 ;
        RECT 4.000 137.000 295.600 138.360 ;
        RECT 4.000 136.360 296.000 137.000 ;
        RECT 4.000 134.960 295.600 136.360 ;
        RECT 4.000 134.320 296.000 134.960 ;
        RECT 4.400 132.920 295.600 134.320 ;
        RECT 4.000 132.280 296.000 132.920 ;
        RECT 4.000 130.880 295.600 132.280 ;
        RECT 4.000 130.240 296.000 130.880 ;
        RECT 4.000 128.880 295.600 130.240 ;
        RECT 4.400 128.840 295.600 128.880 ;
        RECT 4.400 127.520 296.000 128.840 ;
        RECT 4.400 127.480 295.600 127.520 ;
        RECT 4.000 126.120 295.600 127.480 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
        RECT 4.000 125.480 296.000 126.120 ;
        RECT 4.000 124.080 295.600 125.480 ;
        RECT 4.000 123.440 296.000 124.080 ;
        RECT 4.400 122.040 295.600 123.440 ;
        RECT 4.000 121.400 296.000 122.040 ;
        RECT 4.000 120.000 295.600 121.400 ;
        RECT 4.000 119.360 296.000 120.000 ;
<<<<<<< HEAD
        RECT 4.000 118.680 295.600 119.360 ;
        RECT 4.400 117.960 295.600 118.680 ;
        RECT 4.400 117.320 296.000 117.960 ;
        RECT 4.400 117.280 295.600 117.320 ;
        RECT 4.000 115.920 295.600 117.280 ;
        RECT 4.000 115.280 296.000 115.920 ;
        RECT 4.000 113.920 295.600 115.280 ;
        RECT 4.400 113.880 295.600 113.920 ;
        RECT 4.400 113.240 296.000 113.880 ;
        RECT 4.400 112.520 295.600 113.240 ;
        RECT 4.000 111.840 295.600 112.520 ;
        RECT 4.000 111.200 296.000 111.840 ;
        RECT 4.000 109.800 295.600 111.200 ;
        RECT 4.000 109.160 296.000 109.800 ;
        RECT 4.400 107.760 295.600 109.160 ;
        RECT 4.000 107.120 296.000 107.760 ;
        RECT 4.000 105.720 295.600 107.120 ;
        RECT 4.000 105.080 296.000 105.720 ;
        RECT 4.000 104.400 295.600 105.080 ;
        RECT 4.400 103.680 295.600 104.400 ;
        RECT 4.400 103.040 296.000 103.680 ;
        RECT 4.400 103.000 295.600 103.040 ;
        RECT 4.000 101.640 295.600 103.000 ;
        RECT 4.000 100.320 296.000 101.640 ;
        RECT 4.000 99.640 295.600 100.320 ;
        RECT 4.400 98.920 295.600 99.640 ;
        RECT 4.400 98.280 296.000 98.920 ;
        RECT 4.400 98.240 295.600 98.280 ;
        RECT 4.000 96.880 295.600 98.240 ;
        RECT 4.000 96.240 296.000 96.880 ;
        RECT 4.000 94.880 295.600 96.240 ;
        RECT 4.400 94.840 295.600 94.880 ;
        RECT 4.400 94.200 296.000 94.840 ;
        RECT 4.400 93.480 295.600 94.200 ;
        RECT 4.000 92.800 295.600 93.480 ;
        RECT 4.000 92.160 296.000 92.800 ;
        RECT 4.000 90.760 295.600 92.160 ;
        RECT 4.000 90.120 296.000 90.760 ;
        RECT 4.400 88.720 295.600 90.120 ;
        RECT 4.000 88.080 296.000 88.720 ;
        RECT 4.000 86.680 295.600 88.080 ;
        RECT 4.000 86.040 296.000 86.680 ;
        RECT 4.000 84.680 295.600 86.040 ;
        RECT 4.400 84.640 295.600 84.680 ;
        RECT 4.400 84.000 296.000 84.640 ;
        RECT 4.400 83.280 295.600 84.000 ;
        RECT 4.000 82.600 295.600 83.280 ;
        RECT 4.000 81.960 296.000 82.600 ;
        RECT 4.000 80.560 295.600 81.960 ;
        RECT 4.000 79.920 296.000 80.560 ;
        RECT 4.400 78.520 295.600 79.920 ;
        RECT 4.000 77.880 296.000 78.520 ;
        RECT 4.000 76.480 295.600 77.880 ;
        RECT 4.000 75.840 296.000 76.480 ;
        RECT 4.000 75.160 295.600 75.840 ;
        RECT 4.400 74.440 295.600 75.160 ;
        RECT 4.400 73.800 296.000 74.440 ;
        RECT 4.400 73.760 295.600 73.800 ;
        RECT 4.000 72.400 295.600 73.760 ;
        RECT 4.000 71.760 296.000 72.400 ;
        RECT 4.000 70.400 295.600 71.760 ;
        RECT 4.400 70.360 295.600 70.400 ;
        RECT 4.400 69.720 296.000 70.360 ;
        RECT 4.400 69.000 295.600 69.720 ;
        RECT 4.000 68.320 295.600 69.000 ;
        RECT 4.000 67.680 296.000 68.320 ;
        RECT 4.000 66.280 295.600 67.680 ;
        RECT 4.000 65.640 296.000 66.280 ;
        RECT 4.400 64.240 295.600 65.640 ;
        RECT 4.000 63.600 296.000 64.240 ;
        RECT 4.000 62.200 295.600 63.600 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.000 60.880 295.600 61.560 ;
        RECT 4.400 60.160 295.600 60.880 ;
        RECT 4.400 59.520 296.000 60.160 ;
        RECT 4.400 59.480 295.600 59.520 ;
        RECT 4.000 58.120 295.600 59.480 ;
        RECT 4.000 57.480 296.000 58.120 ;
        RECT 4.000 56.120 295.600 57.480 ;
        RECT 4.400 56.080 295.600 56.120 ;
        RECT 4.400 55.440 296.000 56.080 ;
        RECT 4.400 54.720 295.600 55.440 ;
        RECT 4.000 54.040 295.600 54.720 ;
        RECT 4.000 53.400 296.000 54.040 ;
        RECT 4.000 52.000 295.600 53.400 ;
        RECT 4.000 51.360 296.000 52.000 ;
        RECT 4.400 50.680 296.000 51.360 ;
        RECT 4.400 49.960 295.600 50.680 ;
        RECT 4.000 49.280 295.600 49.960 ;
        RECT 4.000 48.640 296.000 49.280 ;
        RECT 4.000 47.240 295.600 48.640 ;
        RECT 4.000 46.600 296.000 47.240 ;
        RECT 4.400 45.200 295.600 46.600 ;
        RECT 4.000 44.560 296.000 45.200 ;
        RECT 4.000 43.160 295.600 44.560 ;
        RECT 4.000 42.520 296.000 43.160 ;
        RECT 4.000 41.160 295.600 42.520 ;
        RECT 4.400 41.120 295.600 41.160 ;
        RECT 4.400 40.480 296.000 41.120 ;
        RECT 4.400 39.760 295.600 40.480 ;
        RECT 4.000 39.080 295.600 39.760 ;
        RECT 4.000 38.440 296.000 39.080 ;
        RECT 4.000 37.040 295.600 38.440 ;
        RECT 4.000 36.400 296.000 37.040 ;
        RECT 4.400 35.000 295.600 36.400 ;
        RECT 4.000 34.360 296.000 35.000 ;
        RECT 4.000 32.960 295.600 34.360 ;
        RECT 4.000 32.320 296.000 32.960 ;
        RECT 4.000 31.640 295.600 32.320 ;
        RECT 4.400 30.920 295.600 31.640 ;
        RECT 4.400 30.280 296.000 30.920 ;
        RECT 4.400 30.240 295.600 30.280 ;
        RECT 4.000 28.880 295.600 30.240 ;
        RECT 4.000 28.240 296.000 28.880 ;
        RECT 4.000 26.880 295.600 28.240 ;
        RECT 4.400 26.840 295.600 26.880 ;
        RECT 4.400 26.200 296.000 26.840 ;
        RECT 4.400 25.480 295.600 26.200 ;
        RECT 4.000 24.800 295.600 25.480 ;
        RECT 4.000 24.160 296.000 24.800 ;
        RECT 4.000 22.760 295.600 24.160 ;
        RECT 4.000 22.120 296.000 22.760 ;
        RECT 4.400 20.720 295.600 22.120 ;
        RECT 4.000 20.080 296.000 20.720 ;
        RECT 4.000 18.680 295.600 20.080 ;
        RECT 4.000 18.040 296.000 18.680 ;
        RECT 4.000 17.360 295.600 18.040 ;
        RECT 4.400 16.640 295.600 17.360 ;
        RECT 4.400 16.000 296.000 16.640 ;
        RECT 4.400 15.960 295.600 16.000 ;
        RECT 4.000 14.600 295.600 15.960 ;
        RECT 4.000 13.960 296.000 14.600 ;
        RECT 4.000 12.600 295.600 13.960 ;
        RECT 4.400 12.560 295.600 12.600 ;
        RECT 4.400 11.920 296.000 12.560 ;
        RECT 4.400 11.200 295.600 11.920 ;
        RECT 4.000 10.520 295.600 11.200 ;
        RECT 4.000 9.880 296.000 10.520 ;
        RECT 4.000 8.480 295.600 9.880 ;
        RECT 4.000 7.840 296.000 8.480 ;
        RECT 4.400 6.440 295.600 7.840 ;
        RECT 4.000 5.800 296.000 6.440 ;
        RECT 4.000 4.400 295.600 5.800 ;
        RECT 4.000 3.760 296.000 4.400 ;
        RECT 4.000 3.080 295.600 3.760 ;
        RECT 4.400 2.360 295.600 3.080 ;
        RECT 4.400 2.215 296.000 2.360 ;
=======
        RECT 4.000 118.000 295.600 119.360 ;
        RECT 4.400 117.960 295.600 118.000 ;
        RECT 4.400 117.320 296.000 117.960 ;
        RECT 4.400 116.600 295.600 117.320 ;
        RECT 4.000 115.920 295.600 116.600 ;
        RECT 4.000 114.600 296.000 115.920 ;
        RECT 4.000 113.200 295.600 114.600 ;
        RECT 4.000 112.560 296.000 113.200 ;
        RECT 4.400 111.160 295.600 112.560 ;
        RECT 4.000 110.520 296.000 111.160 ;
        RECT 4.000 109.120 295.600 110.520 ;
        RECT 4.000 108.480 296.000 109.120 ;
        RECT 4.000 107.120 295.600 108.480 ;
        RECT 4.400 107.080 295.600 107.120 ;
        RECT 4.400 106.440 296.000 107.080 ;
        RECT 4.400 105.720 295.600 106.440 ;
        RECT 4.000 105.040 295.600 105.720 ;
        RECT 4.000 104.400 296.000 105.040 ;
        RECT 4.000 103.000 295.600 104.400 ;
        RECT 4.000 102.360 296.000 103.000 ;
        RECT 4.000 101.680 295.600 102.360 ;
        RECT 4.400 100.960 295.600 101.680 ;
        RECT 4.400 100.280 296.000 100.960 ;
        RECT 4.000 99.640 296.000 100.280 ;
        RECT 4.000 98.240 295.600 99.640 ;
        RECT 4.000 97.600 296.000 98.240 ;
        RECT 4.000 96.240 295.600 97.600 ;
        RECT 4.400 96.200 295.600 96.240 ;
        RECT 4.400 95.560 296.000 96.200 ;
        RECT 4.400 94.840 295.600 95.560 ;
        RECT 4.000 94.160 295.600 94.840 ;
        RECT 4.000 93.520 296.000 94.160 ;
        RECT 4.000 92.120 295.600 93.520 ;
        RECT 4.000 91.480 296.000 92.120 ;
        RECT 4.000 90.800 295.600 91.480 ;
        RECT 4.400 90.080 295.600 90.800 ;
        RECT 4.400 89.440 296.000 90.080 ;
        RECT 4.400 89.400 295.600 89.440 ;
        RECT 4.000 88.040 295.600 89.400 ;
        RECT 4.000 87.400 296.000 88.040 ;
        RECT 4.000 86.000 295.600 87.400 ;
        RECT 4.000 85.360 296.000 86.000 ;
        RECT 4.400 84.680 296.000 85.360 ;
        RECT 4.400 83.960 295.600 84.680 ;
        RECT 4.000 83.280 295.600 83.960 ;
        RECT 4.000 82.640 296.000 83.280 ;
        RECT 4.000 81.240 295.600 82.640 ;
        RECT 4.000 80.600 296.000 81.240 ;
        RECT 4.000 79.920 295.600 80.600 ;
        RECT 4.400 79.200 295.600 79.920 ;
        RECT 4.400 78.560 296.000 79.200 ;
        RECT 4.400 78.520 295.600 78.560 ;
        RECT 4.000 77.160 295.600 78.520 ;
        RECT 4.000 76.520 296.000 77.160 ;
        RECT 4.000 75.120 295.600 76.520 ;
        RECT 4.000 74.480 296.000 75.120 ;
        RECT 4.400 73.080 295.600 74.480 ;
        RECT 4.000 71.760 296.000 73.080 ;
        RECT 4.000 70.360 295.600 71.760 ;
        RECT 4.000 69.720 296.000 70.360 ;
        RECT 4.000 69.040 295.600 69.720 ;
        RECT 4.400 68.320 295.600 69.040 ;
        RECT 4.400 67.680 296.000 68.320 ;
        RECT 4.400 67.640 295.600 67.680 ;
        RECT 4.000 66.280 295.600 67.640 ;
        RECT 4.000 65.640 296.000 66.280 ;
        RECT 4.000 64.240 295.600 65.640 ;
        RECT 4.000 63.600 296.000 64.240 ;
        RECT 4.400 62.200 295.600 63.600 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.000 60.160 295.600 61.560 ;
        RECT 4.000 59.520 296.000 60.160 ;
        RECT 4.000 58.160 295.600 59.520 ;
        RECT 4.400 58.120 295.600 58.160 ;
        RECT 4.400 56.800 296.000 58.120 ;
        RECT 4.400 56.760 295.600 56.800 ;
        RECT 4.000 55.400 295.600 56.760 ;
        RECT 4.000 54.760 296.000 55.400 ;
        RECT 4.000 53.360 295.600 54.760 ;
        RECT 4.000 52.720 296.000 53.360 ;
        RECT 4.400 51.320 295.600 52.720 ;
        RECT 4.000 50.680 296.000 51.320 ;
        RECT 4.000 49.280 295.600 50.680 ;
        RECT 4.000 48.640 296.000 49.280 ;
        RECT 4.000 47.280 295.600 48.640 ;
        RECT 4.400 47.240 295.600 47.280 ;
        RECT 4.400 46.600 296.000 47.240 ;
        RECT 4.400 45.880 295.600 46.600 ;
        RECT 4.000 45.200 295.600 45.880 ;
        RECT 4.000 44.560 296.000 45.200 ;
        RECT 4.000 43.160 295.600 44.560 ;
        RECT 4.000 41.840 296.000 43.160 ;
        RECT 4.400 40.440 295.600 41.840 ;
        RECT 4.000 39.800 296.000 40.440 ;
        RECT 4.000 38.400 295.600 39.800 ;
        RECT 4.000 37.760 296.000 38.400 ;
        RECT 4.000 36.400 295.600 37.760 ;
        RECT 4.400 36.360 295.600 36.400 ;
        RECT 4.400 35.720 296.000 36.360 ;
        RECT 4.400 35.000 295.600 35.720 ;
        RECT 4.000 34.320 295.600 35.000 ;
        RECT 4.000 33.680 296.000 34.320 ;
        RECT 4.000 32.280 295.600 33.680 ;
        RECT 4.000 31.640 296.000 32.280 ;
        RECT 4.000 30.960 295.600 31.640 ;
        RECT 4.400 30.240 295.600 30.960 ;
        RECT 4.400 29.560 296.000 30.240 ;
        RECT 4.000 28.920 296.000 29.560 ;
        RECT 4.000 27.520 295.600 28.920 ;
        RECT 4.000 26.880 296.000 27.520 ;
        RECT 4.000 25.520 295.600 26.880 ;
        RECT 4.400 25.480 295.600 25.520 ;
        RECT 4.400 24.840 296.000 25.480 ;
        RECT 4.400 24.120 295.600 24.840 ;
        RECT 4.000 23.440 295.600 24.120 ;
        RECT 4.000 22.800 296.000 23.440 ;
        RECT 4.000 21.400 295.600 22.800 ;
        RECT 4.000 20.760 296.000 21.400 ;
        RECT 4.000 20.080 295.600 20.760 ;
        RECT 4.400 19.360 295.600 20.080 ;
        RECT 4.400 18.720 296.000 19.360 ;
        RECT 4.400 18.680 295.600 18.720 ;
        RECT 4.000 17.320 295.600 18.680 ;
        RECT 4.000 16.680 296.000 17.320 ;
        RECT 4.000 15.280 295.600 16.680 ;
        RECT 4.000 14.640 296.000 15.280 ;
        RECT 4.400 13.960 296.000 14.640 ;
        RECT 4.400 13.240 295.600 13.960 ;
        RECT 4.000 12.560 295.600 13.240 ;
        RECT 4.000 11.920 296.000 12.560 ;
        RECT 4.000 10.520 295.600 11.920 ;
        RECT 4.000 9.880 296.000 10.520 ;
        RECT 4.000 9.200 295.600 9.880 ;
        RECT 4.400 8.480 295.600 9.200 ;
        RECT 4.400 7.840 296.000 8.480 ;
        RECT 4.400 7.800 295.600 7.840 ;
        RECT 4.000 6.440 295.600 7.800 ;
        RECT 4.000 5.800 296.000 6.440 ;
        RECT 4.000 4.400 295.600 5.800 ;
        RECT 4.000 3.760 296.000 4.400 ;
        RECT 4.400 2.895 295.600 3.760 ;
      LAYER met4 ;
        RECT 23.295 31.455 97.440 269.785 ;
        RECT 99.840 31.455 174.240 269.785 ;
        RECT 176.640 31.455 251.040 269.785 ;
        RECT 253.440 31.455 279.385 269.785 ;
>>>>>>> 5f73601 (Re-hardened with latest Zube version.)
  END
END zube_wrapped_project
END LIBRARY

